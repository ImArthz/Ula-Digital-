-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Oct 18 15:05:40 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY shifter IS 
	PORT
	(
		INPUT :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MIR :  IN  STD_LOGIC_VECTOR(35 DOWNTO 0);
		N :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC;
		OUTPUT :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END shifter;

ARCHITECTURE bdf_type OF shifter IS 

COMPONENT decoder2_4
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 S0 : OUT STD_LOGIC;
		 S2 : OUT STD_LOGIC;
		 S1 : OUT STD_LOGIC;
		 S3 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	OUTPUT_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SLL8_OUT :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SRA1_OUT :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(0 TO 7);


BEGIN 
SYNTHESIZED_WIRE_11 <= "00000000";



OUTPUT_ALTERA_SYNTHESIZED <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


Z <= SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_5;


b2v_inst11 : decoder2_4
PORT MAP(A => MIR(22),
		 B => MIR(23),
		 S0 => SYNTHESIZED_WIRE_10,
		 S2 => SYNTHESIZED_WIRE_6,
		 S1 => SYNTHESIZED_WIRE_7,
		 S3 => SYNTHESIZED_WIRE_9);


SYNTHESIZED_WIRE_2 <= SLL8_OUT AND (SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6);


SYNTHESIZED_WIRE_0 <= SRA1_OUT AND (SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_7);


SYNTHESIZED_WIRE_1 <= INPUT AND (SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8);


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;

SLL8_OUT(31 DOWNTO 8) <= INPUT(23 DOWNTO 0);



SLL8_OUT(7 DOWNTO 0) <= SYNTHESIZED_WIRE_11;



SYNTHESIZED_WIRE_3 <= NOT(OUTPUT_ALTERA_SYNTHESIZED(31) OR OUTPUT_ALTERA_SYNTHESIZED(30) OR OUTPUT_ALTERA_SYNTHESIZED(29) OR OUTPUT_ALTERA_SYNTHESIZED(27) OR OUTPUT_ALTERA_SYNTHESIZED(28) OR OUTPUT_ALTERA_SYNTHESIZED(26) OR OUTPUT_ALTERA_SYNTHESIZED(24) OR OUTPUT_ALTERA_SYNTHESIZED(25) OR OUTPUT_ALTERA_SYNTHESIZED(23) OR OUTPUT_ALTERA_SYNTHESIZED(21) OR OUTPUT_ALTERA_SYNTHESIZED(22) OR OUTPUT_ALTERA_SYNTHESIZED(20));

SRA1_OUT(30 DOWNTO 0) <= INPUT(31 DOWNTO 1);



SYNTHESIZED_WIRE_4 <= NOT(OUTPUT_ALTERA_SYNTHESIZED(19) OR OUTPUT_ALTERA_SYNTHESIZED(18) OR OUTPUT_ALTERA_SYNTHESIZED(17) OR OUTPUT_ALTERA_SYNTHESIZED(15) OR OUTPUT_ALTERA_SYNTHESIZED(16) OR OUTPUT_ALTERA_SYNTHESIZED(14) OR OUTPUT_ALTERA_SYNTHESIZED(12) OR OUTPUT_ALTERA_SYNTHESIZED(13) OR OUTPUT_ALTERA_SYNTHESIZED(11) OR OUTPUT_ALTERA_SYNTHESIZED(9) OR OUTPUT_ALTERA_SYNTHESIZED(10) OR OUTPUT_ALTERA_SYNTHESIZED(8));

SRA1_OUT(31) <= INPUT(31);



SYNTHESIZED_WIRE_5 <= NOT(OUTPUT_ALTERA_SYNTHESIZED(7) OR OUTPUT_ALTERA_SYNTHESIZED(5) OR OUTPUT_ALTERA_SYNTHESIZED(6) OR OUTPUT_ALTERA_SYNTHESIZED(4) OR OUTPUT_ALTERA_SYNTHESIZED(2) OR OUTPUT_ALTERA_SYNTHESIZED(3) OR OUTPUT_ALTERA_SYNTHESIZED(1) OR OUTPUT_ALTERA_SYNTHESIZED(0));

N <= OUTPUT_ALTERA_SYNTHESIZED(31);
OUTPUT <= OUTPUT_ALTERA_SYNTHESIZED;

END bdf_type;